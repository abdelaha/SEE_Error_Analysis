
// n_0
module Cone_n_0 (n_0, i_2_ );
	input i_2_;
	output n_0;
	INVX1 g2088(.IN (i_2_), .QN (n_0));
endmodule

