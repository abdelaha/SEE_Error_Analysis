
// n_3
module Cone_n_3 (n_3, i_3_, i_8_ );
	input i_3_, i_8_;
	output n_3;
	ISOLANDX1 g2084(.ISO (i_3_), .D (i_8_), .Q (n_3));
endmodule

