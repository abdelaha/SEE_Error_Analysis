
// n_4
module Cone_n_4 (n_4, i_5_ );
	input i_5_;
	output n_4;
	INVX2 g2089(.IN (i_5_), .QN (n_4));
endmodule

