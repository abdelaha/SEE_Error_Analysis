
// n_12
module Cone_n_12 (n_12, i_6_ );
	input i_6_;
	output n_12;
	INVX4 g2090(.IN (i_6_), .QN (n_12));
endmodule

