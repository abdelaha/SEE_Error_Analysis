
// n_7
module Cone_n_7 (n_7, i_3_, i_8_, i_0_ );
	input i_3_, i_8_, i_0_;
	output n_7;
	wire n_3;
	NOR2X4 g2082(.IN1 (n_3), .IN2 (i_0_), .QN (n_7));	ISOLANDX1 g2084(.ISO (i_3_), .D (i_8_), .Q (n_3));
endmodule

