
// n_5
module Cone_n_5 (n_5, i_4_, i_7_ );
	input i_4_, i_7_;
	output n_5;
	ISOLANDX2 g2085(.ISO (i_4_), .D (i_7_), .Q (n_5));
endmodule

