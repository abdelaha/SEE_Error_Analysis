
// n_1
module Cone_n_1 (n_1, i_0_, i_5_ );
	input i_0_, i_5_;
	output n_1;
	NAND2X1 g2087(.IN1 (i_0_), .IN2 (i_5_), .QN (n_1));
endmodule

